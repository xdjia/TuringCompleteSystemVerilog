// ComponentFactory
// Is a tool, not a challenge!