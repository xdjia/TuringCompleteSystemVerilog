// The very first level of Turing Complete.

module CrudeAwakening (
    input logic x, output logic y
);
    assign y = x;
endmodule