// Basically a register.

module SavingGracefully (
    input logic clk, save, value,
    output logic outputs
);
    
    DelayedLines register ()
endmodule